� �   �������������������EE�����������������EFEEF���EEEEFFEFEEEEEFFEEFEEEEEEEEEEFEFEEEEEFFE��F����FFFEEE�������������������������������������������������������������EFEEEEFFEFEEEFEEEE������EEEEEEEEFEFFEEFFEEEEEE���������EEEEEF�������FFEFEEFEFEEFFEFFEF�����EEEFE��������������������EE����������������FEEEEF���EEEEFEEFEEEEEFFEEFE��������������F���EE����������F������EFEF���FEEEEFEEEFEEFFFEFFEFFEFFFFFFEFEEEEEEFFEE�������FEEEEE��������������������������������������������������������������FEEEEFEEEFEEEEEE�����E�EFFEEEEEFEEEFFFFEEEF�����������FEEEE��������FEFEEEFFEEFFFEFEEF����EEFFFE����������������F���EE�����������������EFEF���FEFEEEEEEFEEFFFEFFEF��������������EEEEF�������������FE����EEEEEFEFEEFEEEFFEEFEFFEFFFEEFFFFFFEFFEEEEEEFEF��������EFEEEEF�������������������������������������������������������������EEEFEEFFEEEEE����EEEEEEEEEEEEFEEEFEEEEEFE�������������EFF���������FFEEFEEEFFFEEFEEEF����EE��������������������EEEE��F��������F�FFE����EEEEEFEFEEFFFEEFFEFEFEEFFE������F������EEEFFF������������FFFF��FFFEEFEEEEEEEFFEFEFEEEEEFEFFEEFFFFFEEFEEEFEFFEEFF������FEFFEE��������������������������������������������������������������EEEEEEFFEEEE����FFFEEFEFEEEFFEEFFEFEEEEE��������������E�������������EEEEEEEEEFEEEEFEEE�F�E������������F������EEFFF�������������FFF����FFEEEEEEEEEEFFEFEFEEEEEFEF�������������EEE�EFFF�����������EE����FEEEEFEEFEFEEEFFEEEFFEFFEEFEFFEFFEEFEEFFEEEEEEF������EEFFEEF����������������������������������������������������������������FEFEEFEEEE����F�EEFEFE��FEEEEEFEEFEEEEF�������������������������F�EFFEEEEEEFEEEEEEEFEEEFF�����������������FEEFFEEFF�����������EE����FFEEEFEEFEFEEEFFEEEFFEFFFF�����������FFEFEE�F�E�������F��FEF����EEFEEEEEEEEEEEFFEEEFEEFFEEEEFEEFEFEEFFEFEEFFEEFEE���EEFEEEE������������������������������EEE����������������������������������EEFEEEEE������EEEEEE���FEFEEFEFEEEEEF����������������������������EEEEEEEFEE�FEEEFFFFEFF����������������FFEEEE��F�����������FEF����EEFEEFEEEEEEEEFFEEEFEFFEEE�������������EEEFEEEE���������F������FEEEFEEEEEEEEEEFEEEEFEFFEEFFFEFEEEFEFEEFFEFFFEFFFE�FFEEEEFEFF����������������������������FEEEF�������������������������������FFEEFEEEE������EEFFEEF���FEEFEEFFEEEEEFF������FE�����������������FEFEFFFEFFF����EEE�EEF��������������������EEEFEEEE���������F�������EEEFEEEEEEEEEEFEEEFFEEFEFF������������EEEEE�FFFE����������������FFEEEEEEFEFEEEEEFEEEFFEEEEEFEEEEEEFEEEEEFEEFEEFEEFFEEEEFEEF�����������������������������FEEE�������������������������������FEEEEEFEE��������EEEEE�����FEEFEEFEEFEEE������FEEE���������������F��E�FFFFEEE��������FEE�������������������EEEEEEFFFE���������������FEFEEEEEEFEFEEEEEFEEEFFEEEE������������E�EFF��EEEF���������������EFEEEEEEEEFEFEEFEEEFFFEEFEEEEFEFEFEEEEFFEEEEEEEE������EEEEEFF����������������������������EEEE������������������������������EEEFEEEFF�������FEEEFEF�����EEFEEE���E�������EEEEEE����������������E��EEFEEEEF�����������������������������E�EFFF�EEEF���������������EFEEFEEEEEFEFEEFEEEFFFEEFF�������������EEEFEFEEF����������������FEEEFEEEEEEEEFEFFFFEEFEEEFEEEEEEFFFFEEFFFEEEEFFF�������EEEE����������EE�F���������������FEFF��������������������������������EEEEEEE������E�EFEE�F������EEEEFF�����������EFEEEF��������������FE�E�FEFEEFEFF�����������������������������EEEF�FEEF����������������FEFEEEEEEEEFEFEFFFFEEFEEEF��F����������FEF��EEEEF���������������FFFEEEEEEEFFFEFEEFFFEFFEEFFEEEFFEFEEEEFEEEFEF������������������������FEE�����������������EFF��������������������������������EEFFFF����������EE����������EEE�F�����������FFEEE�������������������E�EFEFEFEE���F��������������F����������FEFFFEEEEF���������������EEFEEEEEEEFEFEFEEFFFFFFEEF��EE����������FEF�EEEE���������������FEEEEEFEFEEEFEEEFFFFFFEE���FEEEEEEEEEEEEEEF����������������������������FF���������������������������������������������������F��FF������������������������EEF��������������EEF������������������������FEEEEEF�����������������EE����������FEF�FFEE���������������FEEEEEFEFEEEFEEEFFFFFEEE����FFEE�����������E���FE����������������EFEEEEEFEFEFEEEEFFFEFEE���FEF��FEFEFEEEF�����������������������������EEE�����������������FF������������������������������������������������������������������������������FEF����������������������������FE�����������������FEEE����������EF���FE����������������EFEEEEEFEFEFEEEEFFFEEEE���EEEEE���������FEF����F�������������F�EEEEEEFEFEE��EEEEEEEEEE����������������F�����������������������������F�F���������������������������������������������������������������������������������������������������������������������������������������������������FFEEE���������EFE����F�������������F�EEEEEEFEFEE��EEEEEEEEEE����EEEEE������������F���F�������������EFEEEEEEFEFEF��������EEE����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������EEEEEE������������F�����������������EFEEEEEEFEFEF��������EEE�����FEEEF����������FEE�����������������EFEEEEFEEFF����������������������������������������������������������F�����������������������������������������������������������������������������������������������������������������������������������������������������FEFEEFF����������FEE�����������������EFEEEEFEEEF������������������FEEFFE��������F�EEE���������������F���EEEFFEF��������������������������������������������������F�������������������������FF���������������������������������������������EF�����������������������������������F�����������������������������������������������EEEEEFFFE��������F�EEE���������������F���EEEFEEF�������������������EEEEEEE�������EEFEE�������������������FEEEEEE�������������������������������������������������������������������������������������������������������������������������EEEF����������������������������������������������������������������������������������FEEEFEEEEEE�������EEFEE�������������������FEEFEEE�������������������FEEFEE��������FFFEF�������������������EEEFFEF�����������������������������������������������EEF����F��EE�������������������������������������������������������������FEEEF���������������������������������F���������������������������������FFF���������F�EFFEFEEEFEE��������EFFEF�������������������EEEEE���������������������EFEEEE���������FEEEE����������������FEFFFE�������������������������������������������������EEEEE�FEF�F���������������������������������������������������������������EEEEF���������������������������������F��������������������������������EFEEEEE������EEF�EEEEFEEEE���������FEEE�����������������FEFFFEF���������������������FFEEEF�F�������EEEEF����������������EEF��E���������������EEFE������������������������������EEEEFEEEEFF���������������������������������������������������������������EEF�������������������������������������������������������������������FEEEEEEEE�����EEEFFEEFFEEEF���������EEEE�����������������EEFF�E���������������EEE����EFEEE�����������FEF�����������������F�FEEE��������������FEEFFE���������FEEEF��������������FEEEEFEEEEE����������������������������������������������������������������EEF�����������������������������������������������������������������FEEEEEEFEFFF����EEEEFEEEFEEE�����������FEF�����������������F�FEEE��������������FEFEEE��EFEFF������������EE�����������������FEEEFF��������������FEEFFE����������EEEFFEFEE����������FEFEFEEEEEE�����������������������������������������������������������������������������������������������������������������������������������FEEEEEFFEFF�����EFEEEEEEFEFF������������EE�����������������FEEEFF��������������FEFFFE��EEEE������������F�������������������F�E�F���������������EEEEEEE������EFFFEEEEEEEE���������FFEEEEEEEEE�����������������������������������������������������������������������������������������������������������������������������������EFEFEEEEEEEEF����EEEEFFFEEEE������������F�������������������F�E�����������������EFEEEEE�EEFEF�������������������������������������������������FEEEEEEEE�����FEEFEFFFEFEEE���������EEEEEEEE��F����������������������������������������������������������������������������������������������������������������������������������FEEEEEEEEEEEE����FEEEEFEEEEFEF��������������������������������������������������EEEEEEE��FEEE�������������������������������������������������EFEEEEFEF������EEEEFFEEEEFEE���������EFEEEEF����������������������������������������������������������������������������������F��������������������������������������������������EFEFFFFFEEEEEE�����FFFEEEFFFEE�������������������������������������������������EEEEEEFEF��EEF��������������������������������������������������EFEEEEF��������EEEFFFFEEEEEF������EF�EE����������������������������������������������������������������������������������������F�������������������������������������������������EEFEFEFEEEEEFFFFF��FFFFFEEEFF��������������������������������������������������EFFEEEF����EF����������������������������������������������������E�FFE���������FFEFEFFFEFEF������EEEE�E�������������������������������������������������������������������������������������������������������F�������������������������������FFEEFFEFEEEEFFEEEE�����EEFEEEEE����������������������������������������������������FFFFE�����������������������������������������������������������FFE�����������EEEFEEEEEEFE�FEF��EEEEFEE������������������������������������������������������������������������������������������������������EF�����FEFFE������EF�����������FEEEEEEEFEEEEEEFEE�����EEEEFF�������������������������������������������������������EFEF�������������������������������������������������������������F�����������FEEEEEEEFEFFFE�EE�FEFEEEE�����������������������������������������������������������������������F��������������������������������E���FEFEEEEE���FFEEFF��������FFEEEEEEEEFEEF���EF������EE�����������������������������������������������������������F���������������������������������������������������������������������������FFFFEEF��EE���FFE��EEFEE��������������������������������������������������������������������������������FF����������������������������FEEEEEEE�EEEEE���E�����FEFEEEEEEEEEEEEE������������������������������������������������F�������������������������������������������������������������������������������������������������F�F��FE����E�����EFEFF��FE����������������������������������������������������������������������F��������������������������������������EEEEEEEEFEEEE����������EEFEEFFFEEEFFFEE�����������������������������������������������F��������������������������������F������������������������������������������������������������������EE�����F���FF���FFEEEF�������������������������������������������������������������������������FF�������������������������������������FEEEFEEEEF�FF����������FEFEEFFEFFFEFEFF����������������F����������������������������������������������������������������EF���������������������������������������������������������������EEFF������F������FEEEF�����������������������������������������������������������������������������������������������������������������FFE�����������������������F������EEEFE������������������EE��������������������������������������������������������������������������������������������������������������������������������EFE����E��������FE�������������������������������������������������������������������������������������������������������������������������������������������������FEEEEEFF����������������������������������������������������������������������������������������������������������������������������������������������������FFEFF�F�FFF�����FEEF�����������������������������������������������������������������������������������������������������������������FF�����������������������������FEEEEEFF�����������������������������������������������������������������������������������F����������������������������������������������������������������FE�EFFEEFEFEFFEEEEEE�����������������������������������������tt�����������������������������������������������������EEEEE����������EEEFEEE���������������������������EFFEFF��������������������F��������������������������������������������������������������F�����������������������������������������������������������������FEFEFEFEEEFFEEEFEFE������������������������������������������t�t����������������������������������������������������FFEFFF����������FF�EEEE��������������������������FEEEEFE������������������F���������������������������������������������������������������������������������������������������������������������������������E�EEEFFFEFEEEEFEEEEF���������������������������������������ttt�t������������������������������������������������������FE����������������FFFE��E����������������������FEEEEEEF�����������������������������������������������������������������������������������������������������������������F��������������������������������FEFFFEEFEEFFFEFEEEE��F��������������������������������������ttt��������������������������������������������������������������������������EEEEEEEF��������������������FEEEEFEE����������������������������������������������������������������������������������������������������������������������������������������������������EEEEFEEEEFFEEEEEEF�������������������������������������������tt�������������������������������������������������������������������������FEEEEEEEF���F���������������FEFEEEEE��������������������������������������������������������������������������������������������������������������������������������������������������EEEFEEEEFEFFFFFEEEFE����������������������������������������tt�����������������������������������������������������������������������������EEFEFFF��������������������FFEEEFEF���������������F����������������������������������������������������������������������������������������EEF����F������������������������������������EEEEEFFEFEFFFEEE������������������������������������������t�������������������������������������������������������������������������������F�E������������������������FEF�EE�����������������������������������������EEF������������������������������������������������������������EEEEF������������������������������������������EEEEEEEEEEEEE������������������������������������������������������������������������������������������������������������������������������F������������������������EE�E�����������������������������������������EEEEF���������������������������������������������������������EEEEEEEFF��F�������������������������������������EEEEEEEFEEFE������������FE�����������������������������������������������������������������������������������������������������������������������������������������EE������������������������������������������EEEEFEEEF������������������������������������������������������EEEEFEEEEE�����������������������������������������FEEEFFEFEF�������������EE���������������������������������������������������������������������������������������������F�������������������������������������������FEF����������������������������������������EEEEEEEEEE������������������������������������������������������EFEEEEEEFE��������������������������������������������EEFEEE��������������E��E����������������������������������������������������������������������������������������EEEEEF�����������������������������������������EFF����������������������������������������EFEFEEEEEE������������������������������������������������������EFEEFFEE����������������������������������F�E��������FEEFFFF���������������������������������������������������������������������������������������������������EEF�EEFEEEFE������������������������������������������EE�����������������������������������������EFEEFEEE����������������������������������F�E������������������EEFFF�E�������������������������������������EE������F��FE�������������������������������������������������������������������������������������������t���������EEEEEEEEEEEEFFE�����������������������������������������������������������������������������������EEEFE��EF�����������������������������������EE������������������EEFEEF�����������������������������������������������FE������������������������������������������������������������������������������������������������������EEEFEFFEEEEEEEEF�����������������������������������������������������������������������������������EEFEEF�����������������������������������������������������������EFF�������������������������������������������������EF������������������������������������������������������������������������������������������������������FEEFFFEFFEEEFEE������������������������������������������������������������������������������������EEFF�����������������������������������������������������������FFF������������������������������������������������������������������������������������������������������������t�tt�����������������������������t������������FEEEEFEEEEEEFF�����������������������������������������FE������������������������������������������FF�F�����������������������������������������������������������FEEE�������������������������������������������������������FF�����������������������������������t�tt�����������t��tt������������������������������������������EEEEEFFEEEFEFF�����������������EF����������������������EE�����������������������������������������FFEE���������������������������������������������������������FFEEEEE�������������������������������������������������������F������������������������������������ttt�t���t��t�����ttt�����������������������������t�����������EEEEEFFFFEE������������������F�FE������������������������E��������������������������������������FEEEEEF���������������������������������������������������������EFFEEEF�����������������������������������������������������������������������������������������������t�tttt���������������������������������������������������FEEEFEEEFEE���������������������FFF����������������������EF��������������F�����������������������EFEEEEF���������������������������������������������������������EEEEEEF���������������������������������������������������������������������������������������������������ttt���������������������������������������������������EEEFFFEEEEF������������������FEFEF������������������������������������EE������������������������EEEEEEF��������������������������������������������������������EEEFEEEE���������������������������������������������������������������������������������������������������������������������������������������������������������EEFEEFEEFFE����������������FEFEFEFEE����������������������������������EF�����������������������EEEFEEE��������������������������������������������������F������EEEEEEEEF������������������������������������F�������������������������������������������������������������������������������������������������������������������FFEEEEFEEEFF���������������FEFFFFEEEF���������������������������������F������������������������EEEEEEEF�������������������������������������F����������EEEEEFF�FFEFEEEEF�����������������������������������E�E���������FFFEE�F�������������������������������������������������������������������������������������������������E�FEFFFEEEE���������������EEFEEFFEEEEF�E�������������������������F����������������������EEEEEFF�FFEFEEFEF�����������������������������������E�E��������EEEEFEFEEEEEEEEEFE����������������������������������FEFE���������EEEEEFE��������������������������������������������������������������������������������������������EE���EEEEFFEFEEEE��F���F�����FEEEEFFFEFFEEEE�E��������������F��������EEE��������������������EEEEFEEEEEEEEEEEFE����������������������������������FEFE��������FEEEFEEFFEEFFEEEEEE���������������������������������EFEEEF������EEEEEEFEEF��������������������������������������������������������������F�������������������������FEEEEFFEEEEFFEFEEEFEEFF����F�F�FEFFEEFEEEEEF������������FEEFFEFEFFEE��EFFFEEEF����������������FFEEFEEFFEEFFEEEEEE���������������������������������EFEEEF������FEEEEEEEEEEFEFEEFFF��������������������������������EF�FEE������FFEEEEFFEEE�������������������������������t��������������������������EEFE�����������������������EEEEEEEEEEEEEFEFFFFEEEEF�F������EEFFEEFFFEFEEFF�����������EEEEEEEEFEEEEEEEEEEFEEE�F��������������FFEEFEEEEEEFEFEEFFF��������������������������������EF�FEE��������EEEEEFEFFEFEFFFFFE����������F���������������������EFEFEE�������FEEEFFEEEE�������������������������������������������������������FFEEFFEE���������������������EFEEEEEEEEEEFEFEEEEFEFEEEEF����EFFEFEEEEFEFFFEEF����������FFEEEEFEEEFEFEEEEFE�EE�FEF��������������EEEEEEEEFFEFEFFFFFE��������������������������������EFEFEE�������EEFEFFEEFEEEEFFFFF�������������������������������FEE�EE�F���������EEFEEEE���������������������������������t�����������������������FEEE�EFEF������������������EEEEEEFFFFEEEEEEEEEEEFEFEEFEEE�FEEEEEEFEEFEFFEEE������������FFEEFEFFEFEFEEFEFE����FF�F��������������EFEFFEEFEEEEFFFEF�������������������������������FEE�EE�F�������EFFEEFFEFFFEFFEEFF�������������������������������FEFEFEEF����������FFEE�����������������������������������tt����������������������������EEFE���������������EFEEFEFFFEFEEEEEEEFFFFEEEEEFEEEEFEEEEFFEFEFEEFFEEF�������������EEEE��EEEEEEFEEEF���������������������EFFEEFFEFFFEFFEEEF�������������������������������FEFEFEEF�������FEEFEEEEFEFEEEEEFF������������������������������EFFEE�FF�������������������������������������������������ttt��������������������������FEEEEE����FFF�������FEEEEEEFEEEEEEEEFEEEFEFFEFFEEFEEEEEEEEEEFEFEFEEEEFF�������������FEEFF�FFFEEFEFE�����������������������FEEFEEEEFEFEEEEFEF������������������������������EFFEE�FF�������FEEFEEEEEEEEEEEEFF��������������������������������FEEEFEE�F�F�����F�������������������������������������tttttt���������������������������FFEE���EFFF�������EFEEFFFFEEEFEEEEEEFEEEEEFFFEFEFEFEEEEFFEEEEFFFEFFFEE������������EEF�FEFEEEFFFEFF���������������������FEEFEEEEEEEEEEEEFF��������������������������������FEEEFEE���F���FEFEFFFEEEEFEEEF����������������������������F����FFEEEFEEFFEE���FEEF�������������������������������������ttttt�����������������������������EEEF���FFF������FEEEEFFEEEFFEEEEEEEEEEFFEFFEEEFEEEFEEFEEEEEEFFFFEFEEEEE�������FEEE�FE�EEEEEEE������������������������FEFEFFFEEEEFEEEF��������������������������E������F�EEEFEEFFFE����EEEEEFEEEEEEEFE�����������������������F�FE��EF����EEFEFEFEFEFF�EEEF�����������������������������������ttttt�����������������������������EEEFEFEE�FEE����EFEEEFFEEFEEEEFEEEEFEFEFEEFEEEEEFEEEEFEEEEFEEFFEEEEFEEFFFFF�����EEEEEEEEFEEEEEEE������������������������EEEEEFEEEEEEEFE�����������������������F�FEE�EE����EEFEFEFEFEEF��EEEFFEEEEFEEEF�����������������������FEEFEFEEE��F�FEEFEEFEEEEEEEEEE������������������������������������ttt������������������������������EEEFFEEFF�EEF���EEEFEFEEEFEEFEEEEFFFEFEFFEFEFFEFFEEEEEFEEFFEEFEEEEFEEEEFFE�����EEFFEFEEEFEEEEFF�������������������������EEEFFEEEEFEEEF������������������������EEFEFFEF��F�FEEFEEFEEEEE����FEFFFEEFEEF�������������������������FEFEEEF��FFEEEEEEEFEEEFF�EFE�������������������������������������tt�������������������������������EEFEFFEF���������EEEEEEEEFFFEFFEEEFEEEEFFEEEEEEEEFFFEEEE���EEFFEFEEFEEEFFFE����FEFFF���FEEEEEF��������������������������F�FEFFFEEFEEF�������������������������FEFEEEF����EEEEEEEFEEFFFF���FEEEEEEEEFEE������������������������EEFEEE����F�EEEE�FEEEEEEF�����������������������������������������t������������������������������EEFEEEEE����������EEEEFEEEEEF�������EEEFFEEEFFEEFEF�E�F������FEEEFEEEEFF�EE�F��EFFEEEEE��FEEFF�������������������������F�FFFEEEEEEEEFEE������������������������EEFEEEF��F�EEEEE�FEEEFEEEEEEEEFEEEEEEEFEEF����������������������EEEEEE����FEFEEEF�EFFFEE������������������������������������������������������������������������FEEEEEEE�����������FEEFEEEFFFF�������E�E��EEFEEEEEEEEF������������FEEEEEE�FE����EEEEEEE�F���FFF�����������������������FEEEEEEEFEEEEEEEEEFF����������������������EEEEEE�����EFEEEF�EFEFFEEE������EEFEEEEFEF�������������������FFEEEEEFF����FEFEFF�FF��EFF�����������������������������������������������������������������������EEEFFEEF�������������FEEFFEEFEF��������F��F�EEEEEEEEEEFF������������FFFEE���FF���EEEEEEF�����EFFF���������������������FEFEE������EEFEEEEFEF�������������������FFEEEEEEE����FEFEF��FF��EEFEE������EEEEFFEFE������������������E�E�FEEEEFF�����FEFEFFE�FEEFE�������������������������������������������������������������������������EEF����������������FEFFFEEFFE������FEFFEEEEFFEFFEEEEEEFFEF��������EFEEEEFF�����FEEEEE��EEEFEEEEFEE����������E����FFEEEEEE������EEEEEFEFE������������������E��EEEEEEFF�����FEFEFEF�FEEEFEE�������E����FEF������������������FFFFFFEFEEF�����F��EF�F��EFEE���������������������������������������������������������������������������������������������FEEEE�FEF�����FEEEEEEEEFEEEEEFEEEE�E�����F�E�FFFEEE��������EEEEEEF�EEEEEEEEEEE�������F��EE���F�EFEEE��������E������F������������������FE�FFFEEEEF�����F��EF�F���FEEE����������������������������������EEEF�FEEEEF��������������FFEE�F����������������������������������������������������������������������������������������������EEEFFF���FEEEEEFEEFEFFFEEFFEEEEF����EF�E�FFEEFEEEE�������FEEEF���FFEFEEFFEE������FFFEEEFEFEFFEFEEF��������������������������������EFEEFF�FEEEF��������������FFEE����������������������������������EF�����FEEEE��������������FFFF����������������������������������������������������������������������������������������������FEFEEE�����EEEEFEEEEEEFFEFFFFEFFFF����EEF�FEFEFFEEFF������FFEEEF����EEEFEEFEEE������EEEEEF�E�FEEEEE����������������������������������F�F���FEEEE��������������FFFFF���������������������������������EF�EEE�EEEEF�����������������������������������������������������������������������������������������������������������������FEEEFE����EFEEEEEEFEEFEFFEEEFFEEE���FFF��EEEEFFFE�������F��FFEF������EEEEEEEFEE��FEEEEF��FE���EFF����������������������������������EE�E�E�EEEEF���������������F��EE�������������������������������EEFEEFE�FEEEE����������������������������������������������������������������������������������������������������������������EEFEEEF����EEFFFEFEEEEEFFEEEFFEEEFF��EEE��E�EEEFFE�F������EEEEE�������FFFFE�FFEEE��EFEEF��E����EEFEE�������������������������������EEFEEEE�FEEEE������������������EF�������������������������������EFEEFFEFFEEE����������������������������������������������������������������������������������������������������������������EEEEEEF������FFFFEEEFFEFFFEEEEFEEEFEFFEFEF���FEEFEEE��������EEEE���������������FEFE�FEEEEEF�FF�EEEEEF�������������������������������EFEEFEEFFEEE�������������������FEE����������������������������FEEEEEEE���FEF����������������������������������������������������������������������������������������������������������������FEFFFEEE�����EEEFFEEFEFEFFEEFFFFEEEFEEEEE�����FEEEEE���������FE����������������EEFEFEEEEEE�F�FFFEFEEEE����������������������������FEFFEEEE���E�F�������������������EFF��������������������������FEEEF�EEEF����������������������������������������������������������������������������������������������������������������������EFEEEEEE�����EFEFEEEEFFEEEFFEFEEFFEEEEFE���������EFEFEE������E����������������EEFEEFEEFFFE�FFEEEEEEFFF��������������������������FEEEF��EEF�������������������������FEEE��������������������������EEEEEEEE���������������������������������������������������������������������������������������������������������������������FFEEFEEFEFFFF��FFEFEFFFFFEFEEEFEFEEEEEEEEFF������������FE������F������������F��FEEEEF�EEE�EFFEEEEEEFEFEE���������������������������EEEEEEEE��������������������������EEE�������������������������FEEEEEEEEEE�������������������������������������������������������������������������������������������������������������������FEEEEFEEEF����FFFEEFEEFEFEEFEEEFEFEEEEEEEEF����������������������������������EEFEEEEEF��F��FFFEEEEFFEEEFF�������������������������FEEEEEEEEEF�������������������������EEFF�����������������������FEEEFEFEE�F�������������������������FFF������������������������������������������������������������������������������FF�������FEEEFFEFEFE���EEEEEEEEFFFEEEEEFEEFEEFEEEEE�E���������������������������������EEEFFEEEEEF�����FEFEEEEEFFEEFF������������������������EEEFEEEEEF������������������������FEFEE������������������������EEEEEEFEE��������������������������EEE��������������������������������������������������������������������������F���FEFEF�����FEEEFFEEFEF��FFEEFEEEFFFFEEEEEEFEEEFFEEFEEFE���������������������������������EEEEEEFEFF�������FFFFFEEFEFEE������������������������EEEEEEFEE��������������������������FEEEE������������������������EEEEEEFFF��������������������������EEEEF�����������������������������������������������������������������������FEFEEFFEEEEFEE�FFEEFFFEEEE��FFFEEEFEFEEEEEE��EFEEEEEFEEE��F����������������������������������EFEEEEEEFF���������EEEEEFEFE�����������������������FEEEEEEFFE��������������������������EEEEEE����������������������FEEEEFFEE���������������������������F�E����������������������������������������������������������������������F�EEEFEEFEEEEEEEEEEEEEFFEEEEFF��EEFEEFEEEFEFE�����FEEFFFEEEE������������������������������������EFEEEEFEEE��������FFEEFEEEEEE����������������������FEEEEFEFF����������������������������FE�������������������������EEEEEEEF�����������������������������FE���������������������������������������������������������������������EEFEEEEFFFEEEEEEEEFEEEFEEEEFFEE��EEEFEFFEFFEEF������EEEEFEEE���������������������������������������EEFE�EF�����������F�EEEEF������������������������EEEEEEEF�����������������������������F��������������������������E��EEFEF���������������������������������������������������������������������������������������������������EEEEFEEFFEFFEFEFEEFEFEEFEEEFEFEF�FEEFFFEFEFFEEEEE����EEEFEE��������������������������������������������������������������E���������������������������F��EEFEF���������������������������������������������������������E����F����������������������������������������������������������������������������������������������������FEEEEEEEEFFFEFFEEFFEEEFFEEEEEEF���EEFEEFEFEFEFEEF����EEEEF���������������������������������������������������������������������������������������������F���F������������������������������������������������������������F��F���������������������������������������������������������������������������������������������������EEEEFEEEEEFEEEEEEEFEEEEFFFEEEFEE���EEEFFEFEEFEEFEEEF��E�F������������������������������������������������������������������������������������������������F��F�������������������������������������������������������������������������������������������������������������������������������������������������������������������EEEEFFFFEEEFEFEFEEEFEFEEEFEEFEEF���FEEEFFFEFEEEFFEEEF���������������t�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������FEEFFFEFEEEEFEFF���EEEEFEEFFFEEF���EEFEFEEFFEEEFEEEEE��������������t������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������EEEFEEEFEFFFEE������FFEEEEEEEEEE��FEEEEEEEFEFEEFFEEEF�������������ttt�����������������������������������������������������������������������������������������������������������������������������������������������������EE����������������������������������������������������������������������������������������������������EEEEFEEEEFEEF��������FEEEEEEEEEFFEEEEEEEEEEEEEEEEEEEF��������������tt�������������������������������������������������������������������������������������FE�������������������������������������������������������������EEE����������������������������������������������������������������������������������������������������FEEEFFFFEFE�����������FFFFEEEEEFEEFEEFFEEFFEEEEEFFEFF�������������t�����������������������EE�������������������������������������������������������������EEE�������������������������������������������������������������EEEF���������������������������������������������������������������������������������������������������FEEEEFEFFFF�������������FFFEEF���EFEEEEEEFEFEEFEEEE���������������������������������������FF�������������������������������������������������������������EEEF�������������������������������������������������������������FEF����������������������������������������������������������������F���������������������������������FEFFEEEFEE����������������FF�������F�FEEFFEEEEE�FF����������������������������������������F�F��������������������������������������������������������������EEF������������������������������������������������������������FEF���������������������������������������������������������������������������������������������������FEFFFEFFFEF�����������FEEFEEEF�������EFEEEFEEEFFF������������������t��������������������FEEEEEF�����������������������������������������������������������FF��������������������������������������������������������������E�F�������������������������������������������������������������������������������������������������FEEFEEFFEFEEEE����������FEEFFEEE������FEEF�FEEEEE��������������������t�������������������F�FEEEEF�����������������������������������������������������������EEF�������������������������������������������������������������EEE�����������������������������������������������F������������������E�������F���������������������EFEEFFFFFEEEE�E�������FF��FFEFEEEE�����F�F��EFEFFFFE����������������������������������������EFEEEF�����������������������������������������������������������EEE���������������������������������������������������������E��FEEE���������������������������������������������������������������������������F�������������������EEEEEEEFFEEEF��EE���F�EFFFFEF��EFEFEF���FF�FEEEEEEEE������������������������������������������FEE���������������������������������������������������������E��FEEE�������������������������������������������������������FEFEE�F�������������������������������������������������������������������������������������������������EEEEEEEEEEF����E����EFEEEFFFE��FE��F����FFFFEFEEEEEF������������������������������������E���������������������������������������������������������������FEFEE�F��������������������������������������������������������EEEEFEEFE�������������������������������������������������������������������������������������������������F�FEFEEEE�����F���FEEEEEEEEEE�FE�FFF��EEEEEEFFFFEE������������������������������������EEF�������������������������������������������������������������EEEEFF�FE�������������������������������������������������������FFEEFEEEE�����������������������������������������������������������������������������������������������������F�EEF���������FEEEEEEEEFEEEFFFFFEFEEEEEEFEFEEF�����������������������������������EEF��������������������������������������������������������������FFEEFEEEEF�����������������������������������������������������EFEEEEEEEEF�����������������������������������������������������������������������������������������������������������������EEEEFEFFFEFFEEEEEEEEEFFFEEEFEEEEF�����������������������������������EEF�������������������������������������������������������������EFEEEEEEEEF��������������������������������F��������������������EEEEFEEFEEE����������������������������������������������������������������������������������������������������������������EEEEEEFEEFEEEEEFFEEEFEFEFFFEFFEEEE�����������������������������������EEF����������������������EF���������������F���������������������EEEEFEEFEEE����������������������������������������������������FEEFFFFEFFE�F���������������������������������������������������������������������������������������������������������������EFEEEEEEFEFFEEEEFEEEFEEEEEEEEEEFFE����������������������������������EEEF������������������EEE�EFF��������������E��������������������FEEFFFFEFFE�F���������������������������������������������������EEFEEEFFFEEFEF�����������������������������������������������������������������������������������������������������������������FEEEFEEEEFFFFFFFFFFEFFFEEEFE�E����������������������������������FEEEF�������������������EEFE������������������������������������FEEFEEEFFFEEFEF������������������������������������������������FEEEEFEFEEEFEEEE������������������������������������������������������������������������������������������������������������������EEEEEEEEEFFFFFFFFEEEFEEFF�������������������������������������EEEEEE������������������FEEFE������������������������������������FFEEFFFEEEFEEEE������������������������������������������������EFEEFEEFEEEFEFEE������������������������������������������������������������������������������������������������������������������FFEEFFEEEFFFEFEEEEFEEEEF��������������������������������������FFFEEFEF�����������������FF�������������������������������������EFEEFEEFEEEFEEFE������������������������������������������������FEFEEEFEEFFEEFF��������������������������������������������������������������������������������������������������������������EEFFEEEF�EEEEEFFFFEEEEEFEFEEE���������������������������������F�FFEEEEEEFEE��������������������������������������������������������FEFEEEFEEFFEEFFE���������������������������������������������������EEEEFEE��FF�F�����������������������������������������������������������������������������������������������������F������FEEEEEEFEEEEEEEEFFFEEEFEEEF�����������������������������������FFFEEEEEEEFFEE�����������������������������������������������������������EEEEFEE��FF������������������������������������������������������EEFEF������������������������������������������������������������������������������������������������������������������EEEEEEEEEEFEEFEEEEFEEEF����������������������������������������FEEEEEEEEEEEE�������������������������������������������������������������EEEEF������������������������������������������������������������FEFE������������������������������������������������������������������������������������������������������������������EEEEEEEEEFFFEFEFEFEEE������������������������������������������FEEEEFFEEEFF���������������������������������������������������������������FEFF������������������������������������������������������������FEEF�������������������������������������������������������������������������������������������������������������������EFEEFEEEEEEEEEEEEEE�������������������������������������������EEEFFEEE�������������������������������������������������������������������FEE��������F��������������������������������������������������FEFFEE���EEEEEF���������������������������������������������������������������������������������������������������������FFEEFEFEEEEEFEEEEE�F������������������������������������������EEEEEFEFF������������������������������������������������������������������EFFEEFF�EEFEEF�������������������������������������������������FEEEEEEEEEEEEEE��������������������������������������������������������������������������������������������������������FEFEEEEEEEEEEEFFFF���������������������������������������������EEEE�FEEF�����������������������������������������������������������������FEEEEEEEEEEEEEE���������������������������������������F�������FEEEFFEEEEFFEEEEF�����������������������������������������������������������������������������������������������������FEEEEFEEEEEEFFFFFEEEF��������������������������������������������EEEEEEE�����������������������EF���������������������������������F�������FEEEFFFEEEFFEEEEF�������������������������������������FEEF����FFEEEEEFFFEEFEFEEE�������������������������������������������������������������������������������������������������������FEFEEEFFFEEEFF��������������������������������������������������EEEEFF�����������������������FEE�������������������������������FEEF�����FFEEEEFFFEEFEFEEEE�������������������������������������EEEFE�F��EFEFEEEEEEEEEEEE�������������������������������������������������������������������������������������������������������F��FEEFEFEEEFEE����������������������������������������������������EFE������������������������EEEE������������������������������EEEFF�F�EEFFEEFEEEEEEEEEEF���������������������������������F��EEEEEEFEEEEEEEEEEFEEEEFEEE����������������������������������������������������������������������������������������������������������FEEFEEEEFEFF�����������������������������������������������������EEF������������������������EFEF�������������������������F��EEEEEEFFEEEEEEEEEEEEEEFEEE���������������������������������EEEFEFFEEEFFEEEEFEEFFEEEFFF�������������������������������������������������������������������������������������������������������������F����FEEEF��������������������������������������������������������FF������������������������FFEEF�����������������������EEEFEFFEEEFFEEEEFEEFFEEEFFF�����������������������������������FFEEEFEEEEFFEEEEEEEFEEEEEEEFEE����������������������������������������������������������������������������������������������������������������EFFF�����������������������������������������������������������F������������������������EFEEF��������������������FFFEEEFEEEEFFEEEEEEEFFEFEEEEFEE����������������������������������EFEFFEEEFEEEFEEEEEEEFFFFEEEEFEE����������������������t�t���������������������������������������������������������������������������������������E�����������������������������������������������������������������������������������FEEEFEEFE������������������EEEFEFFEEEFEEEFEFEEEEEEFFFEEEEFEE����������������������ttt��������EFEFFFFEEEFEEFEFFFFEFEFEEEEEFF������������������������t����������������������������������������������������������������������������������������������������������������������������������������������F����������������������������EEEEEEEEEE����������������EEEEEFEFFFFEEEFEEFEFFFFEEEFEEEEEFF������������������������t���������FEEEEFFFEFFEEEFEEFEEEEEEEEFEEE��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������FF�E�FEFEFEEE�F�����������FEEFEEFEEEEFFFEFFEEEFEEFEEFEEEEEFEEE����������������������������������EFEFFFFFFEFFFEEFEFEEFFFFEEEEE���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������FEFEEFFEEEEEEFF�����������EEEEFFEFEFFFFFFEFFFEEFEFEEFFFFEFEEE�����������������������������������FEFFFFFFFEFFEFFEEEFFFEEEEEFE������������������������������������������������������������������������������������������������������������������������������������FF��E�F����������������������������������������������������������F�EEE�FFEEFEEFFF�����EFEFEEEEEEFEFFFFFFFEFFEEFEEEFFFEEEEEF�������������������������������������FEFFFFEEEFFEEE�FFFEEFFEEEEF���������������������������������������������������������������������������������������������������������������������������������F��EFEFFEEEFEF�FFE������������������������������������������������������FEF�EEFFEEF�������FEEEFEEFEEEEFFFFEEEFFEEE�FFFEEFFFEEEF�������������������������������������FFFFEEEFEE�E���������FEFE�����������������������������������������������������������������������������������������������������������������������FF����������EFEEEEEEEFEEFEFEFEEEE��������������������������������������������������������EFFEF��������EEEEFEEEFFFFFFEEEFEE�E��������FFEEE���������������������������������������EFFEFEF���������������FF���������������������������������������������������������������������������������������������������������������������FEFEEFE�EEEEEEEEEFEEEEEEEEEEEFEEEEEEEE���������������������������������������������������������F�����������EEFFEEFFEFFEFEF����������������F����������������������������������������EEEEEE���������������������������������������������������������������������������������������������������������������������������������������FEEEEEEEEEEEFEEEEFEEFFEEEEEEEEFFEEEEEE������������������������������������������������������������������������FEEEEEEEEEE����������������������������������������������������������EEEEEF���������������������������������������������������������������������������������������������������������������������������������������FFEEEEEEEEEEFEEFEFEFEEEEEEEEFFFFFEFEFEF������������������������������������������������������������������������EEEFEEFEFF����������������������������������������������������������EEEEE���������F���������������������������������������������������������������������������������������������������������������������������������EEEEEEEFEFFFFFEFFEEFEEEEEFFEFFFEEEEF������������������������������������������������������������������������FFEEEEEEE�����������������������������������������������������������FFEFE������������������������������������������������������tt��������������������������������������������������������FFF��������������������FE��FFEFEEEEFFFEFEEEEEEFEEEEFFEFFEFEEF���������������������������������������������EE�������������������������FFEFEEFFEFE��������F���������������������������������������������tt���EEEF��������E���������������������������������������������t�tt������������������������������������������������������FFF���������������������F�F�FEFEEFFEEEEEEEFEEFFFFEFEEFEEFEEFE���������������������������������������������FEEE�F������������������EE�FEEEEEEEEEE��������E���������������������������������������������t�tt��EEFF��������F�����������������������������������������t�tt����t������������������������������������������������������FF����������������������F�EEEEFFEEFEFEEEEEFEFFEEEEFEEEEEFFE����������������������������������������������EEEEF��������������������EFEEEEFEEEEFF����������������������������������������������������tt����t�EEEF������������������������������������������������t�ttt��������������������������������������������������EFEEE���FEF������������������������EEEEEFFEFEFFEEFEEEE��EEEEFE�EF���������������������������������������������������FFEEF���EEEFE���������FFEEEFEEEEEEEEF�������������������������������������������������tttt�������FEE��������������������������������������������������tttt������������������������������������������������EEEEEEEF�FE�EF����������������������FFFEEEEEFFFFEEFEFEEE��FF�F��F�������������t��������������������������������������FEEEEE��FFFEEEFEEEF��FEEEEEEEEFEEEFEE��������������������������������������������������t�tt�������EEE��������������������������������������������������ttt��������������������������������������������������EEEEEE����EE����������������������FFFFEEEEFFEEFFEEFEEEFF��������������������t���������������������������������������EEEE����EEEFEEEFEEEE��EEEEEFEFEEEEEEE��������������������������������������������������ttt��������FFF�������E�F���������������������������������������������������������������������������������������������FEEEFE����E�����������������������EEFFFFFFEEEFFFFFEFEEEEF����FE�������������tt��������������������������������������E�EE����FEEEEEEFEEEEE�EEEEEFEEEEEEEFF��������E�������������������������������������������t��������EFEE�����EE�FFF�������������������������������������������������������������������������������������������FFFFE�������E��������������������FEFEEFEEEEEEEEEEEFEFEEFFFEEF��������������t��������������������������FE������������EEFEFF���FEEEFEEEFEEEEEEEEEEFFEEFFEFEE�����EE�FFF�������������������������������������������������EEEE����EEFEE����������������������������������������������������������������������������������������������EEEEF�����������������������EFFF�EEEEEEFFFFEEEFFFEEFFFE��EEEEFF������������������������������������EFEEF������������EEEEE���EEEEE��FFFEEFFEFFEFEFEEEFEFEE����FEEEE���������������������������������������������������FEEEEEFEEEEEEE���������������������������������������������������������������������������������������������EFFF������������������������EEFF�EFEEEEFEEEEEEEFFEF���EEF�F�FFF��������������������������������������EE������F������FEEFF����FEEF�����EEEE���EEFEEEFEEEEF�EFEEEEEEE��������������������������������������������������FEFFEEEFEEEEE���������������������������������������������������������������������������������������������FEEFEE������������������������EE��EFEEEFEEEEEEEFEEE�EFEEF�FEE����������������������������������������EEF������FFE���FEFF�F��FEEFE������FEEF���EEEEFFFEEEEFFEEEEEEEE���������������������������������������������������FFFF��E�EFEEF�����������������������������������������������������������������������������������������FF���EFFEEE�EF��������������������FE��EFEFF�FEEEEEEFEEEEEEFEEFE���������������������������������������������������FEEEEEFEEF����EEEE������FFFEFFF�EFEEEFEEFFEFE�E�EFEEF���������������������������������������������������EFEEF��F�FE���������������������������������������������������������������������������������������FEE�E���EEFEEFEEE���������������������������EFEEFFEEEEEFEFF�EEEEEF����������������������������������������������������FFFEEFFEEE����FEE��������FEE�EFFEEFFFEEEEFEF�����FE�����������������������������������������������������FEEF�����������������������������������������������������������������������������������F�F��������FEEEE���EEEEEFFEEF���������������������������EEE��FEEEEEEE��FFEEE����������������������������������������������������F�EEFEEFFEEE����F��������FEFFEEEEFEEEEEFFFEEE������������������������������������������������������������FEEF����������������������������������������������������������������������������������F�EFF�������EEEEE����FEEEFEEF����������������������������F�F����FEEFFF��F�������������������������������������������������������EE�EEEEF�FFEEEF���F������FEFEEEFFEEEEEEFFFEEEE������������������������������������������������������������EEE������������������������������������������������������������������������������������EEEE������EEEEEE����EFEEFF�E�������������������������������������������F�����������������������������������������������������������EF��FEEEE������������EEEFEEFFFFFEEFFFEEFF�������������������������������������������������������������EE������������������������������������������������������������������������������������FEEFEF������EFEFF���FFEEEEEEE����������������������������������������F���������������������������������������������������������������FF��EFEFF����������FEEEEEEFFEFFEEEEFEEE��������������������������������������������������������������E�������������������������������������������������������������������������������������EFEEEEEF��EFF�����������EFFEE�����������������������������������������������������������������������������������������������������������EEFFF����������FEEFEFEEEEE���EEEEEEF��������������������������������������������������������������EF����������������������������������������������������������������������������������FEEEFFF�F�FE�EF��������������F�����������������������������������F����������������������������������������������������EE�������FFE�������FEFF�����������FFEEEEFEEEF����FFEEEEF��������������������������������������������������������������������������������������������������������������������������������������������������EEEEFE�FFEEEFFF������������������������������������������������FFEF�F������������������������������������������������EEEE�F�EEFFEE�������F��������������FEEEEEEEEEE�FFEFEF������������������������������������������������������������������������������������������������������������������������������������������������������EEEFEE��FFEE��F������������������������������������������������FFF�F���������������������������������������������E��EEFEFEEEEEFFE����������������������EEFFEFEFE����FFEE����������������������������������������������������������������������������������������������������������������������������������������������������F���FEEFFEF���EEEFE���������������������������������������������F�EEE�����������������������������������������������E���EEEEFEEEEEFEE���������������������EEEF�EEEEEF����FEEF������������������������������������������������������������������������������������������������������������������������������������������������EEFFFFFEEEEFF��FFFE��F���F���������������������������E������������FFFEEEF�����F����������������������������������������EFE�FFFEEEEF�FEE������������������������FE�EEF���������F������������������������������������������������������������������������������������������������������������������������������������������������FEEEEEFEEEEE���FFFEEEEE������FEE��������������������EF�����������EEEEFFEEE�������F��������������������������������������FEEE���FFEF������������������������������F�������������������������������������������������������������������������������������������������������������������������������������������������������������FEEEEFEEEEEEE��FEEFEEFFF�����F��E���������������������E�������EFF��EEEEEEEFE�����E����������������EF��������������������EEEE����FEEF�����������������������������������������������������������������������������������������������������������������������������������������������������������������������F������������������EEEEFEFFEEEEFEEFFFEEEEEEFEF���FFFF��������������������������������E��EEFE��FE�����FEEE������������������������������������EEEEE������E�F�����������������������������������������������������������������������������������������������������F��������������������������������������������������������������FF����������������FFFFEFEEEEFEEEEEFEFFEEFEEFEFEFFFEE������������������F�������������������������������EEFE�����������������������������������EEEEFF�������������������������������������������������������������������������������������������������������������FF�����������������������������������������������������������FEEEE���������������FFEEFEEEEEEEEEEEFF����EEEEEEEEEEFF����������������EE�F�������������������������������EEEFF�������������F���������������������EFEEEE�������������������������������������EE������������������������������������������������������������������FEEEE�����������������������������������������������������������FEFF��������������FEEEEEFFFEEFFEFEEE������FEEEEEEFFEE�F������������FEEEEEF�������������������������������FEEEE��������������E������������������FFEEEEE������������������������������������EFFEFF����������������������������������������������������������������FEFFF��������������������������������������������������������FEEFEFE��������������FFEEEFFFEFFFFEFEEF������EEEFEEEFFEE��������������FEEEFF�F�������������������������������FEEE�������������EEE������������������FEFEFEE�����������������������������������FFEEEEFE������������������������������������������������������������EEFEF��F�������������������������������������������������������EEEFE����������������FEFEEFFFEFFFFEEFF��������EEF��EFFE����������������EFEEF��������������������������������EEEEF�������������EFE�����������������FEEEFEFE����������������������������������FEEEEFEEE�����������������������������������������������������������EEEFEF����������������������������������������������������������EEEEF�����������������EFFEFEEEEEEEEFEE�������FF���FF�������������������EEEEE��������������������������������EEEEE�������������EEE������������EE�F�FEFFFFFF�����������������������������F����EEEEEEFE�������������F����������������������������������������������EEEEF�����������������������������������������������������������EEEE������������������FEEEEEEEFEEFEEE�������������FEEE����������������EEEEE�������������F����������F�������EEEEEFF�����EE�FF���EE������������EEFF�FEF�����F�������������������������FEEEEFFFEFFFEEE������������FF�����������������������������������������������EEEE������������������������������������������������������������F����������������������EEF�E�EFEEEEFF��������������EF����������������EFEEF����������EFF�F����������EEF��EFEFEEEEEF�����EEFEF���F���������EFEEFEE�E�EEEE���������������F��������������EEEEEEFEFFEEEF�������������F�����������������������������������������������F����������������������������������������������������������������F��������������������������������F��������������FEFEE���������������FEEE����������EEFF�����������EFEEEFEEEEEEFFEF���F�EEEEEF�����������E�FEEEEFE�EEEEF���������������E��������������EEEEEEEEEEEEE���������������������������������������������������������������F���������������������������������������������������������������E����������������������E��F�F�F���������������EEEEFEEE��������������FEE�F���������FEFFF����������EEEFEEEEEFEEEEEEF��EEE�FE�����F����������FFEEFEE����F��������������FF�����������E�FEEEEFFFEFEEE���������������������������������������������������������������FE��������������������������������������������������������������FE����������������������F���E�E��������������EEEEEEFFEE��������������EEEF����������FEEEF��������F�EEFEEEEEEFFEFFEE����F���E����������������EEEEFEFF��F�������������������������EEEEEFEEEEFEFFEEF����������������������������������������������������������������FFF�����������������������������������������������������������������������������������EEF����F�������������FEFEFFFEEFEF���������������E�F����������FEEEE���������EEEFEEFFEFFFFFEEEE��FFEE������������������EFFEEEF����������������������������EEEEEEFFFFFEEEFFE��������������������������������������������������������������������������������������������������������������������������������������������������������E������F�����������FEEFEEFEEFEEE��������������F�FF����������EEEEF�������FEEEEEEEFFFEFFFEEEEF���FEF�F����������������FEEEEF����������������������������FEEEFEFFFFFFEEEFEE����������������������������������������������������������������������������������������������������������������������������������������������������EEEEE������������������FE�EEEEEFFEEEFF�������������EFEE���������EEEFF�������F�EEEEEEEEFFEFEFEFFF������������������������FFEFEE����������������������������FEEFEEFFFFFEEFEFE���������������������������������������������������������������������������������������������������������������������������������������������������FEFFEEFF�����F������������FEFEEEEEEFEEFF�������������EFE����������FFEEE��������FEFFEEEEEEEFEEEEE������E�����F�������������EFFFEEF�������������������������F�FEEFEEFEFFEEFEFFFF��������������������������������������������������������������������������������������������������������������������������������������������������FEFEFEEE�������EFF�FFF����FF��EEEEEFEEEF���������������������������EFE����������FFFEFEEEFEEEEFEEEF��������F���������������FEEEEE�������������������������FFFFEFFFFFFFFEFEEF�F���������������������������������������������������������������������������������������������������������������������������������������������������EEFEEFEE�����EFEEEEFFFFEEEEE��FEEEEEEEF������������������������������������������F�EEEFFEEEFE�EEEF�����F��F��������������FEFEEF��������E�����������������FFEEFEEEEEEEEEEEF�������������������������������������������������������������������������������������������������������������������������������������������������������FEEFFF������EEEFEEEEEEEEEEEEF�EFEFEEF�������������������������������������������FF�F�EFFFFE�EFEEF�����EEEE�������������FEEFEEEF������F�������������������EEEEEFEFFEEEEF���������������������������������������������������������������������������������������������������������������������������������������������������������FEE��F����FEEEEFEEEEEEFEEEFFFFEFEFEF���������������������������������������������E��������E�EFEEF����FEEEE�������������EEEEEEE��������FF������������������FFEEEEEF�E�F��������������t��������������������������������������������������������������������������������������������������������tt��������������������������������EEEE�������EEEEEEEEEEF�EFEEE�FEEEEEFE�����������������E���������������������������E����F�FEFFFEEEF�F��EFEEF�������������EEFEEEEF�����������������������������EEEEEEEEF��������������tt����������������������������������������tt�������������������������������F������������������������������t���������������������������������EEEF������FFEFEFEEF����EFFFFFEEFEEEEF�������������F�F��F�������������������������FEEFFEEEEEEEFFEEEE���FFEE��������������FEEEEEEEF����������������������������FEFFEEEFF��������������tt����������������������������������������t�������������������������������������������������������������������������������������������������EFEE������������E������FEFF���F�EEF��������������FFE�FF�������������������������EFEEFFFEEEEEFEEEEEE���EEEE��������������EEEFEEEFF������������������������������FFE�F������������������������������������������������������������������������������������������������������������������������������������������������������������EFF������������������������������E���������������EEE���������������������������EEEEEEFEEFEFEEEEEEFF����EFE��������������EFEEEEE�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������E�������������������EFF��������������������������F��FE���������������EF����������������������������EEEEEEEEEEEEFEEEEF������������������������EFFEEF���������������������������������������������������������������������������������������������������������������F����������������F���������������������������������������E�EEEFFE�����������������FE����������������������������������������������FEE����������������������������EEEEEFFFFEEEFFEEE�������������������������EEEFE������������������������������F��������������������������������������������������������������������������FEEEEFF�����������������������EEE����������������������������FEEFFFEEEEEE����������������E�����������������������������������������������������������������������������FFEEFFEEEFFEEEEFE��������������������������EEEE���������������������������FFEEE�EEFE���������F���������������EEF�������EEE����������������������������FEFEFEEEEEEE������������������FFEEEEF���������������������������EEFFFEEEEEEE���������������E�F��������������������E�������������������������E��������������������������F��FEEEEFEEEFEEEEEFF���������������������������EEE�������������������������EEFEEEF�EEFE��������E�F��������������FFE����FFEEEEFF��������������������������EEFFFEEEFEEE���������������E��EEFFFEFEEF������������������������EEFEEFEEEEEEE�������������EFEEE�������������������EEE�����������������������F����������������������������EEEFEEEEEEEFEEEEEE��������������������������F�F��������������������������EFEEE���E�E��������FEFEF��������������F�FF��EEFFFEFEEF������������������������EEEEEEEEEEEEE�������������EF�EEEEEFFFEEF�����������������������FEEEEEEEEEEFEE�������������FEEEE��������������������EE���������������������������������������������������FEFEEEEEEEEFEEFEEEF��������������������������������������������������������FEFF�������������EEEEE���������������FEEE�FEEEEFFEEEF�����������������������FEEFEEEEEEEFEE�������������FE�EEEEEEFFEEE�����������������������FEEFEFEEEEFF�������������FFEEEE�������������������FF��F�������������������������������������������������F�EFEEEEEEEEEEEEEFF���������������������������������������������������������������������������EEE�����������������EEEE�EEEEFFEEEE�����������������������FEEFEFEEEEFF�������������FFEEFEFFFFFFFFEE�����������������������FFFEFEFFEFF�������F�����FEEFEEE�������������������FF��������������������������������������F�F�������������EFEEEEEFEEEEEEFFF���������������������������������������������������������������������������F��������������������E�FEEEFFEEEFFE�����������������������FFEEFEFEEFE��������������EEEE�FFFEFEEEEEF�����������������������F�EFEFEEEEEF�������������EFFEE�������������������FE�������������������������������������������������������EFFFEEEEFEFEEEE�����������������������������������������������������������������������������������������������������FFFEFEEEEEF�����������������������F�EEEFEEEEEF�������������EEFEFFEEFFFFE���������������������������EEFFFFEEEEFFE�����������EEFEE����������������������������������������������������������������������������EEEEFE�������������������������������������������������������������������������������������������������������������FFEEFFFFE���������������������������EEFFFFEEFF�FE����������FEEFEEFEFFEFEE���������������������������EEEFEEEEFF��F������������EEEE���������������������������������������������������������F������������������E��EF������������������������������������������������������������������������������������������������������������F�EFEFFEFEE���������������������������EEEFEEEEFF��F������������EEEFFFFFFE�E����������������������������EEEFEEFFF�FF������������EFF�����������������������������������������������������������F�����������������EF�����������������������������������������������������������������������������������������������������������F�F�FEFFEFFFE�E����������������������������EEEFEEFFF�FE������������EFEFEFFEFFEEF��������������������������FEEFFFEF��FEE������������E�E���������������������������������������������������������F������������������EFF����������������������������������������������������������������������������������������������������������FF�EEEEFEFFEFFEEF��������������������������FEEFFFF����FEF����������EFF�EFFEEEEEFFE�������������������������FFEFEFFF����F������������F�E���������������������������������������������������������F������������������������������������������������������������������������������������������������������������������������������E�FFFEFEEFFEEEEEFFE�������������������������FFEFEFFF����F������������F�E